`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/22/2022 04:21:37 PM
// Design Name: 
// Module Name: zero_counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module varzcount #(parameter WIDTH = 64) (
    input [WIDTH-1:0] hash,
    output [$clog2(WIDTH):0] num_zeros
    );
    
    integer c;
    integer i;
    always @(*) begin: counter
        c = WIDTH;
        i = 0;

        for(i = 0; i < WIDTH; i = i + 1) begin
            if(hash[WIDTH - 1 - i]) begin
                c = i;
                disable counter;
            end
        end
    end
    
    assign num_zeros = c[$clog2(WIDTH):0];
    
endmodule

module zero_counter #(parameter BLOCK_SIZE = 64)(
    input [255:0] hash,
    
    output reg [31:0] num_zeros
    );
    
    // In order to do this more efficiently, we break up our
    // computation into four blocks, and then combine them appropriately.
    // Hopefully, this leads to a more balanced implementation than
    // naively generated by the compiler.
    
    // Create zero counters for four segments of this hash
    wire [$clog2(BLOCK_SIZE):0] counts [256 / BLOCK_SIZE - 1 : 0];
    
    genvar i;
    generate
        for(i = 0; i < 256 / BLOCK_SIZE; i = i + 1)
            varzcount #(BLOCK_SIZE) counter (hash[i*BLOCK_SIZE +: BLOCK_SIZE], counts[i]);
    endgenerate
    
    integer j;
    always @(*) begin: counter
        num_zeros = 32'd256;
        for(j = 0; j < 256 / BLOCK_SIZE; j = j + 1) begin
            if(!counts[(256 / BLOCK_SIZE) - j - 1][$clog2(BLOCK_SIZE)]) begin
                num_zeros = {23'b0,
                             j[7 - $clog2(BLOCK_SIZE) : 0],
                             counts[(256 / BLOCK_SIZE) - j - 1][$clog2(BLOCK_SIZE) - 1 : 0]};
                disable counter;
            end
        end
    end
    
endmodule
